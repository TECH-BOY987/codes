# KERNEL: start reset
# KERNEL: done resetting
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=154    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=77    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=236    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=73    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: rd_en=1    dout=0    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: rd_en=1    dout=0    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=248    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=227    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=57    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______GENERATOR_______
# KERNEL: --------------
# KERNEL: rd_en=1    dout=0    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=154    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=154    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=154    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=77    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=77    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=77    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=236    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=236    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=236    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=73    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=73    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=73    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=154    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=154    empty=0
# KERNEL: --------------
# KERNEL: Scoreboard: Expected Data = 154, Received Data = 154
# KERNEL: Scoreboard: Test Passed for Data = 154
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=154    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=77    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=77    empty=0
# KERNEL: --------------
# KERNEL: Scoreboard: Expected Data = 77, Received Data = 77
# KERNEL: Scoreboard: Test Passed for Data = 77
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=77    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=248    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=248    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=248    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=227    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=227    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=227    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=57    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=57    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: wr_en=1    d_in=57    full=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: ________DRIVER________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=236    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=236    empty=0
# KERNEL: --------------
# KERNEL: Scoreboard: Expected Data = 236, Received Data = 236
# KERNEL: Scoreboard: Test Passed for Data = 236
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=236    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=73    empty=0
# KERNEL: --------------
# KERNEL: Scoreboard: Expected Data = 73, Received Data = 73
# KERNEL: Scoreboard: Test Passed for Data = 73
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=73    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=248    empty=0
# KERNEL: --------------
# KERNEL: Scoreboard: Expected Data = 248, Received Data = 248
# KERNEL: Scoreboard: Test Passed for Data = 248
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=248    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=227    empty=0
# KERNEL: --------------
# KERNEL: Scoreboard: Expected Data = 227, Received Data = 227
# KERNEL: Scoreboard: Test Passed for Data = 227
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=227    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=0
# KERNEL: --------------
# KERNEL: Scoreboard: Expected Data = 57, Received Data = 57
# KERNEL: Scoreboard: Test Passed for Data = 57
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=0
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: Scoreboard: FIFO is empty, no data to read
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: Scoreboard: FIFO is empty, no data to read
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: Scoreboard: FIFO is empty, no data to read
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: Scoreboard: FIFO is empty, no data to read
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: --------------
# KERNEL: _______monitor__________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# KERNEL: Scoreboard: FIFO is empty, no data to read
# KERNEL: --------------
# KERNEL: _________scoreboard___________
# KERNEL: --------------
# KERNEL: rd_en=1    dout=57    empty=1
# KERNEL: --------------
# RUNTIME: Info: RUNTIME_0068 $finish called.