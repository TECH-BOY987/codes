// Code your testbench here
// or browse Examples
`include "uvm_macros.svh"
import uvm_pkg::*;
module tb;
initial begin
  `uvm_info("tb_top","hello world",UVM_MEDIUM);
end
endmodule

"""output"""

# KERNEL: UVM_INFO /home/runner/testbench.sv(7) @ 0: reporter [tb_top] hello world 
