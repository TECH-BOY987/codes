module example;
string s1="HELLO WORLD";
initial begin
    $display("display string s1:%0s",s1);
end
endmodule
